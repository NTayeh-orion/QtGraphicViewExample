module sync_debouncer (input clk, rst_n, input btn_raw, output reg btn_debounced); reg [19:0] counter; reg last_btn; always @(posedge clk or negedge rst_n) if (!rst_n) begin counter <= 0; last_btn <= 0; btn_debounced <= 0; end else begin if (last_btn != btn_raw) counter <= 0; else if (counter < 20d999_999) counter <= counter + 1; else btn_debounced <= btn_raw; last_btn <= btn_raw; end endmodule
