module sync_ram #(parameter ADDR_WIDTH=8, DATA_WIDTH=16) (input clk, input we, input [ADDR_WIDTH-1:0] addr, input [DATA_WIDTH-1:0] din, output reg [DATA_WIDTH-1:0] dout); reg [DATA_WIDTH-1:0] mem [0:(2**ADDR_WIDTH)-1]; always @(posedge clk) if (we) mem[addr] <= din; always @(posedge clk) dout <= mem[addr]; endmodule
