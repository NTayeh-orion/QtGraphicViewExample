module sync_fifo #(parameter DATA_WIDTH=8, DEPTH=16) (input clk, rst_n, input [DATA_WIDTH-1:0] din, input wr_en, rd_en, output [DATA_WIDTH-1:0] dout, output full, empty); reg [DATA_WIDTH-1:0] mem [0:DEPTH-1]; reg [$clog2(DEPTH):0] wr_ptr, rd_ptr; wire wr_full = (wr_ptr == {~rd_ptr[$clog2(DEPTH)], rd_ptr[$clog2(DEPTH)-1:0]}); wire rd_empty = (rd_ptr == wr_ptr); assign full = wr_full; assign empty = rd_empty; always @(posedge clk or negedge rst_n) if (!rst_n) wr_ptr <= 0; else if (wr_en && !wr_full) begin mem[wr_ptr[$clog2(DEPTH)-1:0]] <= din; wr_ptr <= wr_ptr + 1; end always @(posedge clk or negedge rst_n) if (!rst_n) rd_ptr <= 0; else if (rd_en && !rd_empty) rd_ptr <= rd_ptr + 1; assign dout = mem[rd_ptr[$clog2(DEPTH)-1:0]]; endmodule
