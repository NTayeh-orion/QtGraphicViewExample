module and3_gate(input x, input y, input g, output z);
    assign z = x & y;
endmodule