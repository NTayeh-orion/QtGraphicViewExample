module sync_divider #(parameter WIDTH=32) (input clk, rst_n, input start, input [WIDTH-1:0] dividend, divisor, output reg [WIDTH-1:0] quotient, remainder, output reg done); reg [WIDTH-1:0] r, q; reg [4:0] count; always @(posedge clk or negedge rst_n) if (!rst_n) begin quotient <= 0; remainder <= 0; done <= 0; count <= 0; end else if (start) begin r <= dividend; q <= 0; count <= WIDTH; done <= 0; end else if (count > 0) begin if (r >= {1b0, divisor}) begin r <= r - divisor; q <= {q[WIDTH-2:0], 1b1}; end else q <= {q[WIDTH-2:0], 1b0}; r <= {r[WIDTH-2:0], 1b0}; count <= count - 1; end else begin quotient <= q; remainder <= r; done <= 1; end endmodule
