module sync_uart_tx #(parameter CLK_FREQ=50_000_000, BAUD=115200) (input clk, rst_n, input tx_start, input [7:0] data_in, output reg tx, output reg tx_done); localparam BIT_TICKS = CLK_FREQ / BAUD; reg [15:0] bit_timer; reg [3:0] bit_idx; reg [8:0] shift_reg; reg busy; always @(posedge clk or negedge rst_n) if (!rst_n) begin tx <= 1; tx_done <= 0; busy <= 0; bit_timer <= 0; bit_idx <= 0; end else if (!busy && tx_start) begin busy <= 1; shift_reg <= {1b0, data_in, 1b1}; bit_idx <= 0; tx_done <= 0; end else if (busy) begin if (bit_timer == 0) begin if (bit_idx < 9) begin tx <= shift_reg[0]; shift_reg <= {1b1, shift_reg[8:1]}; bit_idx <= bit_idx + 1; bit_timer <= BIT_TICKS - 1; end else begin busy <= 0; tx_done <= 1; tx <= 1; end end else bit_timer <= bit_timer - 1; end endmodule
