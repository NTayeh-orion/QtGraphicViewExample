module add(input [3:0] a, input [3:0] b, input x , input y , input z , output [4:0] sum , output flag , output zer_f , output m);
    assign sum = a + b;
endmodule