module jtag_interface (
    input tck,
    tms,
    tdi,
    output reg tdo,
    input trst_n
);  // IEEE 1149.1 JTAG TAP controller interface
endmodule
