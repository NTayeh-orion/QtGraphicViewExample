module sync_multiplier #(parameter WIDTH=16) (input clk, rst_n, input [WIDTH-1:0] a, b, input start, output reg [2*WIDTH-1:0] product, output reg done); reg [3:0] state; parameter IDLE=0, CALC=1, FINISH=2; always @(posedge clk or negedge rst_n) if (!rst_n) begin state <= IDLE; product <= 0; done <= 0; end else case (state) IDLE: if (start) begin state <= CALC; done <= 0; end CALC: begin product <= a * b; state <= FINISH; end FINISH: begin done <= 1; state <= IDLE; end endcase endmodule
