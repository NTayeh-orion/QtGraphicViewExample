module sync_fsm_moore (input clk, rst_n, input a, b, output reg y); parameter S0=2b00, S1=2b01, S2=2b10, S3=2b11; reg [1:0] state, next_state; always @(posedge clk or negedge rst_n) if (!rst_n) state <= S0; else state <= next_state; always @(*) case (state) S0: next_state = a ? S1 : S0; S1: next_state = b ? S2 : S0; S2: next_state = a ? S3 : S0; S3: next_state = b ? S0 : S3; default: next_state = S0; endcase always @(*) case (state) S0: y = 0; S1: y = 0; S2: y = 1; S3: y = 1; default: y = 0; endcase endmodule
